library verilog;
use verilog.vl_types.all;
entity executeTOmem_sv_unit is
end executeTOmem_sv_unit;
