library verilog;
use verilog.vl_types.all;
entity memoryTOwrite_sv_unit is
end memoryTOwrite_sv_unit;
