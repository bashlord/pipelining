library verilog;
use verilog.vl_types.all;
entity fetchTOdecode_sv_unit is
end fetchTOdecode_sv_unit;
