library verilog;
use verilog.vl_types.all;
entity decodeTOexecute_sv_unit is
end decodeTOexecute_sv_unit;
